/*
   Hazard Unit
*/

module hazard_unit(
    input CLK, nRST,
    hazard_unit_if.hif
);


endmodule
