/*
  Pat Sabpisal
  ssabpisa@purdue.edu
*/

`ifndef PCIFVH
`define PCIFVH

`include "cpu_types_pkg.vh"

interface pc_if;

  import cpu_types_pkg::*;

endinterface

`endif
