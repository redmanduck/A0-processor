/*

  Pat Sabpisal
  ssabpisa@purdue.edu

*/
`include "datapath_cache_if.vh"
`include "cpu_types_pkg.vh"

module control_unit (
   input CLK, nRST,
   datapath_cache_if.cache dcif
);

   import cpu_types_pkg::*;

endmodule
